module main

import cpu

fn main() {
	c := cpu.Cpu.new()
	println(c)
}

module main

import cpu

fn main() {
	println('Hello World!')
}
